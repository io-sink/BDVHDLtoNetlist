library IEEE;
use IEEE.std_logic_1164.all; 

entity 7425ic is 
port (
	attribute library_name : string;
	attribute component_name : string;
	attribute footprint_name : string;
	attribute const_assign : string;
	attribute pin_assign : integer;

	attribute library_name of 7425ic is "74xx";
	attribute component_name of 7425ic is "74HC25";
	attribute footprint_name of 7425ic is "Package_DIP:DIP-14_W7.62mm_Socket_LongPads";

	GND : in std_logic;
	attribute const_assign of GND is "GND";
	attribute pin_assign of GND is 7;
	VCC : in std_logic;
	attribute const_assign of VCC is "VCC";
	attribute pin_assign of VCC is 14;

	1G : in std_logic;
	attribute const_assign of 1G is "VCC";
	attribute pin_assign of 1G is 3;
	2G : in std_logic;
	attribute const_assign of 1G is "VCC";
	attribute pin_assign of 1G is 11;

	1A : in std_logic;
	attribute pin_assign of 1A is 1;
	1B : in std_logic;
	attribute pin_assign of 1B is 2;
	1C : in std_logic;
	attribute pin_assign of 1C is 4;
	1D : in std_logic;
	attribute pin_assign of 1D is 5;
	1Y : out std_logic;
	attribute pin_assign of 1Y is 6;

	2A : in std_logic;
	attribute pin_assign of 2A is 9;
	2B : in std_logic;
	attribute pin_assign of 2B is 10;
	2C : in std_logic;
	attribute pin_assign of 2C is 12;
	2D : in std_logic;
	attribute pin_assign of 2D is 13;
	2Y : out std_logic;
	attribute pin_assign of 2Y is 8
	);
	end 7425ic;

architecture logic of 7425ic is 
begin 

	1Y <= not(1A or 1B or 1C or 1D);
	2Y <= not(2A or 2B or 2C or 2D);

end logic;